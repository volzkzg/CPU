`timescale 1ns/1ps

module test();
    reg clock, reset;

   min_sopc sopc(
        .clk(clock),
        .rst(reset)
    );

    always #1 clock = ~clock;

    initial begin
        $dumpfile("dump.vcd");

        $dumpvars;
       /*
        $dumpvars(0, sopc.cpu.register.storage[1]);
        $dumpvars(0, sopc.cpu.register.storage[2]);
        $dumpvars(0, sopc.cpu.register.storage[3]);
        $dumpvars(0, sopc.cpu.register.storage[4]);
        */
        $readmemh("rom.txt", sopc.inst_rom0.inst_mem);

        clock = 1'b0;
        reset = 1'b1;

        #20 reset = 1'b0;
        #12 `AR(1, 32'h00008000); `AR(2, 32'hxxxxxxxx); `AR(3, 32'hxxxxxxxx); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000000); `AR(2, 32'hxxxxxxxx); `AR(3, 32'hxxxxxxxx); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'hxxxxxxxx); `AR(3, 32'hxxxxxxxx); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h00008000); `AR(3, 32'hxxxxxxxx); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000000); `AR(3, 32'hxxxxxxxx); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'hxxxxxxxx); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h00000000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h00000011); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h00000000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h00000000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h80000010); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h0000000F); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h00000011); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'h00000000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h80000010); `AR(2, 32'h80000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h0000FFFF); `AR(2, 32'h80000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h80000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h00000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h00000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h00000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h00000000); `AR(2, 32'h00000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h00000000); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h00000000); `AR(2, 32'h00000020); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h00000020); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFF); `AR(2, 32'h00000020); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFF); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFF); `AR(2, 32'h00000020); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hA1000000); `AR(2, 32'h00000020); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hA1000000); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hA1000000); `AR(2, 32'h00000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h11000000); `AR(2, 32'h00000001); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h11000000); `AR(2, 32'h00000003); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h11000000); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'h0000FFFF); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFF0000); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFB); `AR(2, 32'h00000000); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFB); `AR(2, 32'h00000006); `AR(3, 32'hFFFF8000); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFB); `AR(2, 32'h00000006); `AR(3, 32'hFFFFFFE2); `AHI(32'h00000000); `ALO(32'h00000000);
        #2  `AR(1, 32'hFFFFFFFB); `AR(2, 32'h00000006); `AR(3, 32'hFFFFFFE2); `AHI(32'hFFFFFFFF); `ALO(32'hFFFFFFE2);
        #2  `AR(1, 32'hFFFFFFFB); `AR(2, 32'h00000006); `AR(3, 32'hFFFFFFE2); `AHI(32'h00000005); `ALO(32'hFFFFFFE2);
        `PASS;
    end
endmodule
